entity test1 is
	port (
		a: in std_logic;
		b: out std_logic_vector(1 downto 0);
		c: out std_logic
		HAHAHAHAHA
	);
end test1;


