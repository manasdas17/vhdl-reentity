library blalalalo.ieee;
use hahaha.ieee;

--tatata tata

entity test2 is
	generic(
		number: integer:=8);
	port (
		--tititi
		c: in std_logic;
		d: out std_logic_vector(3 downto 0)
	); --foo bar
end entity;

architecture foo of test2 is
begin
end architecture;

--tatata

