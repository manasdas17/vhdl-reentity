entity test1 is
	port (
		a: in std_logic;
		b: out std_logic_vector(1 downto 0)
	);
end test1;


